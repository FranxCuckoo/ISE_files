----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:47:19 11/20/2015 
-- Design Name: 
-- Module Name:    oqpsk - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: O-QPSK with halfsine pulse shaping.
--						To form the offset between I-phase and Q-phase chip modulation, the Q-phase
--						chips shall be delayed by Tc with respect to the I-phase chips
--		Combined oqpsk_clocked_v2.vhd and sine.vhd from vhdl examples folder
--		For calculation of sine values: i)  t=0 : pi/10 : 2*pi array of 20 values of time.
--										ii) int32(sin(t) * 127) take the int values
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.trans_pkg.all;

entity oqpsk is
    Port (clk_2Mhz	: in STD_LOGIC;
		  clk_1Mhz	: in STD_LOGIC;
		  reset		: in STD_LOGIC;
		  chip_in	: in  STD_LOGIC;
		  modulation_en : in std_logic;
		  
   		  stream_out : out std_logic 
	
		);
end oqpsk;

architecture Behavioral of oqpsk is
	-- Declaring in-module signals
	signal buffer_iq : STD_LOGIC_VECTOR(1 DOWNTO 0);
	signal en_iq_out : std_logic := '0' ;
	
	-- Number of clk_2Mhz_period to delay
	constant Delay : integer := 1;
	signal delay_buffer_chip : std_logic_vector(Delay downto 0);
	signal quadrature_delayed : std_logic;

	-- Sin and cos signals
	constant clk_sincos_period : time := 0.05 us;
	
	signal clk_sincos : std_logic;
	signal inphase	:  STD_LOGIC;
	signal quadrature : STD_LOGIC;
	signal sine : integer range -128 to 127;
	signal cos  : integer range -128 to 127;
	signal modul_i : integer range -128 to 127;
	signal modul_q : integer range -128 to 127;

	type memory_type is array (0 to 38) of integer range -128 to 127; 
	type memory_type2 is array (0 to 38) of integer range -128 to 127; 
	
	-- ROM for storing the sine values generated by MATLAB. 21 values
	signal pos_sine_values : memory_type := (0, 20, 39, 58, 75, 90, 103, 113, 121, 125, 127, 125, 121, 113, 103, 90, 75, 58, 39, 20, 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);
	signal neg_sine_values : memory_type := (0,-20,-39,-58,-75,-90,-103,-113,-121,-125,-127,-125,-121,-113,-103,-90,-75,-58,-39,-20,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

	signal sine_values : int32_vector (0 to 38) := (0,39,75,103,121,127,121,103,75,39,0,-39,-75,-103,-121,-127,-121,-103,-75,-39,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);
	signal cos_values : int32_vector (0 to 38) := (127,121,103,75,39,0,-39,-75,-103,-121,-127,-121,-103,-75,-39,0,39,75,103,121,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);
	
	-- Convolution signals
	signal modul_q_array : int32_vector (0 to 38) := (others => 0);
	signal modul_i_array : int32_vector (0 to 38) := (others => 0);
	signal convolution_q : int32_vector (0 to 38) := (others => 0); -- (modul_q_array'length + sine_values'length - 2));--38
	signal convolution_i : int32_vector (0 to 38) := (others => 0);
	signal sum : int32_vector (0 to 38) := (others => 0);

begin
	--------------------------------------
	-- Clock process for sinusodials
	--------------------------------------
	clk_sincos_process : process
	begin
	 	clk_sincos <= '1';
	 	wait for clk_sincos_period/2;
	 	clk_sincos <= '0';
	 	wait for clk_sincos_period/2;
	end process;
	
	--------------------------------------
	-- generation of I,Q signals
	--------------------------------------
	INPUT_CHIPS: process(clk_2Mhz)
		variable pointer : integer := 0;
	begin
		if rising_edge(clk_2Mhz) then
			if reset = '1' then
				en_iq_out <=  '0';
				buffer_iq <= "00";
				pointer := 0;
			else
				-- Holding two chips
				buffer_iq(pointer) <= chip_in;

				if pointer = 0 then
					pointer := pointer + 1;
					en_iq_out <= '0';
				elsif pointer = 1 then
					en_iq_out <= '1';
					pointer := 0;
				end if;
			end if;

		end if;
	end process;
	
	OUTPUT_SIGNALS: process(clk_1Mhz, en_iq_out, buffer_iq)
	begin
		if rising_edge(clk_1Mhz) then
			if reset = '1' then
				inphase <=  '0';
				quadrature <= '0';
			else
				-- Output signals for multiplication with sin,cos
				if en_iq_out = '1' then
				 	inphase <= buffer_iq(0);
				 	quadrature <= buffer_iq(1);
				end if;
			end if;
		end if;
	end process;
	
	--------------------------------------
	-- generation of a Tc delay
	--------------------------------------
	delay_buffer_chip(0) <= quadrature;

	gen_delay_en: for i in 1 to Delay generate
		delay_chip: process(clk_2Mhz)
			begin
				if rising_edge(clk_2Mhz) then
					delay_buffer_chip(i) <= delay_buffer_chip(i-1);
				end if;
			end process;
	end generate;

	quadrature_delayed <= delay_buffer_chip(Delay);

	--------------------------------------
	-- Multiplication of sine and chip
	-- Half-pulse shaping of chip data
	-- MSK filtering
	--------------------------------------
	HALF_SIN_MODU: process(clk_sincos)
		variable j : integer range 0 to 20;
		variable w : integer range 0 to 20;
		variable h : integer range 0 to 20;
		variable y : integer range 0 to 20;
	begin
		-- Each rise, outputting a point of sine
		-- we output 20 values out of 21. 
		-- in sin it works due to the common point (0)
		-- but in cos we output 127, ..., 121. We are missing a value,
		-- we should output 127, ..., 127
		if rising_edge(clk_sincos) then
			if reset = '1' then
				modul_i <= 0;
				modul_q <= 0;
				j := 1;
				w := 20;
				h := 1;
				y := 20;
			else
				-- if I want to use sine as a carrier just change 10 to 20.
				case inphase is
				   when '0' => 
					  -- ouputting 10 values.
					  -- 1-10 index
					  modul_i <= neg_sine_values(w);
					  if (w = 1) then
					      w := 20;
					  else
					      w := w - 1;
					  end if;

				   when others => 
					  -- ouputting 10 values.
					  -- 10-1 index
					  modul_i <= pos_sine_values(j);
					  if (j = 20) then
						  j := 1;
					  else
						  j := j + 1;
					  end if;
					  
			    end case;
	
				case quadrature is
				-- If we use cos: Look when signal changes state (1->0, 0->1)
				-- you have mistep, from 127 to -121 and from -127 to 121.
				-- because we dont have the commmon sample as in sin, the 0.
				   when '0' => 
					  -- Different LUT when signal is 0
					  modul_q <= neg_sine_values(y);
					  if (y = 1) then
					      y := 20;
					  else
					      y := y - 1;
					  end if;

				   when others => 
					  modul_q <= pos_sine_values(h);

					  if (h = 20) then
						  h := 1;
					  else
						  h := h + 1;
					  end if;
					  
			    end case;
				
		   end if;
				
		end if;
	end process;

	--------------------------------------------------
	-- Convolution of modulated inphase and modulated
	-- quadrature phase signals. Every 2Tc have an output
	--------------------------------------------------
	Convolving_signals : process(clk_sincos)
	begin
		if rising_edge(clk_sincos) then
			if reset = '1' then
				convolution_q <= (others => 0);
				convolution_i <= (others => 0);
			-- outputting when 127 so the convolution start not at
			-- the beginning of the cos but at the middle(Tc delay)
			elsif (modul_q = 127) or (modul_q = -127) then
				convolution_q <= conv(modul_q_array,sine_values);
				convolution_i <= conv(modul_i_array,cos_values);
			end if;
		end if;
	end process;

	----------------------------------------------------------------
	-- Getting quadrature array of modul_q and modul_i
	----------------------------------------------------------------
	modul_q_array(0) <= modul_q;
	modul_i_array(0) <= modul_i;

	gen_modululated_array : for i in 1 to 19 generate
		process(clk_sincos)
		begin
			if rising_edge(clk_sincos) then
				modul_q_array(i) <= modul_q_array(i-1);
				modul_i_array(i) <= modul_i_array(i-1);
			end if;
		end process;
	end generate;

	--------------------------------------------------
	-- Addition of the two modulated signals
	-- the .* in matlab. point to point multiplication
	--------------------------------------------------
	SUMMING_MOD_SIGS : for j in 0 to 38 generate
	   process(clk_sincos)
	   begin
		   if rising_edge(clk_sincos) then
			   if reset = '1' then
				   sum(j) <= 0;
	   		   else
				-- should connect to stream_out
   				   sum(j) <= convolution_i(j) + convolution_q(j);
			   end if;
		   end if;
	   end process;
    end generate;
	
	----------------------------------------------------------------
	-- TX_enable_delayed = modulation_en
	-- We delayed it again by 8us until the mudul_i and q are ready
	----------------------------------------------------------------
--	delay_modulation_en(0) <= modulation_en;
--
--	gen_delay_chip: for i in 1 to 80 generate
--		delay_chip: process(clk_sincos)
--		begin
--			if rising_edge(clk_sincos) then
--				delay_modulation_en(i) <= delay_modulation_en(i-1);
--			end if;
--		end process;
--	end generate;
--	convolution_en <= delay_modulation_en(80);

	--------------------------------------
	-- generation of sine&cos signals
	-- (not needed really - just for me)
	--------------------------------------
--	GEN_SINE: process(clk_sincos)
--		variable i : integer range 0 to 20 := 0;
--	begin
--		-- Each rise out a point of sine
--		if rising_edge(clk_sincos) then
--			if reset = '1' then
--				sine <= 0;
--				cos <= 0;
--				i := 0;
--			else
--				sine <= sine_values(i);
--				cos <= cos_values(i);
--				i := i + 1;
--				
--				if(i = 20) then
--					i := 0;
--				end if;
--			end if;
--		end if;
--	end process;

end Behavioral;

