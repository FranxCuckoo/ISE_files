----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:47:19 11/20/2015 
-- Design Name: 
-- Module Name:    oqpsk - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: O-QPSK with halfsine pulse shaping.
--						To form the offset between I-phase and Q-phase chip modulation, the Q-phase
--						chips shall be delayed by Tc with respect to the I-phase chips
--		Combined oqpsk_clocked_v2.vhd and sine.vhd from vhdl examples folder
--		For calculation of sine values: i)  t=0 : pi/10 : 2*pi array of 20 values of time.
--										ii) int32(sin(t) * 127) take the int values
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity oqpsk is
    Port (clk_2Mhz	: in STD_LOGIC;
		  clk_1Mhz	: in STD_LOGIC;
		  reset		: in STD_LOGIC;
		  chip_in	: in  STD_LOGIC;
		  modulation_en : in std_logic;
		  
   		  stream_out : out std_logic	
	
		);
end oqpsk;

architecture Behavioral of oqpsk is
	-- Declaring in-module signals
	signal buffer_iq : STD_LOGIC_VECTOR(1 DOWNTO 0);
	signal en_iq_out : std_logic := '0' ;
	
	-- Number of clk_2Mhz_period to delay
	constant Delay : integer := 1;
	signal delay_buffer_chip : std_logic_vector(Delay downto 0);
	signal quadrature_delayed : std_logic;

	-- Sin and cos signals
	constant clk_sincos_period : time := 0.10 us;
	
	signal clk_sincos : std_logic;
	signal inphase	:  STD_LOGIC;
	signal quadrature : STD_LOGIC;
	signal sine : integer range -128 to 127;
	signal cos  : integer range -128 to 127;
	signal modul_i : integer range -128 to 127;
	signal modul_q : integer range -128 to 127;

	type memory_type is array (0 to 10) of integer range -128 to 127; 
	
	signal sum : integer range -256 to 255;
	
	-- ROM for storing the sine values generated by MATLAB. 21 values
	signal pos_sine_values : memory_type := (0,39,75,103,121,127,121,103,75,39,0);
	signal neg_sine_values : memory_type := (0,-39,-75,-103,-121,-127,-121,-103,-75,-39,0);
	-- signal cos_values : memory_type := (127,121,103,75,39,0,-39,-75,-103,-121,-127,-121,-103,-75,-39,0,39,75,103,121,127);
	-- signal inv_cos_values : memory_type := (-127,-121,-103,-75,-39,0,39,75,103,121,127,121,103,75,39,0,-39,-75,-103,-121,-127);

begin
	--------------------------------------
	-- Clock process for sinusodials
	--------------------------------------
	clk_sincos_process : process
	begin
	 	clk_sincos <= '1';
	 	wait for clk_sincos_period/2;
	 	clk_sincos <= '0';
	 	wait for clk_sincos_period/2;
	end process;
	
	--------------------------------------
	-- generation of I,Q signals
	--------------------------------------
	INPUT_CHIPS: process(clk_2Mhz)
		variable pointer : integer := 0;
	begin
		if rising_edge(clk_2Mhz) then
			if reset = '1' then
				en_iq_out <=  '0';
				buffer_iq <= "00";
				pointer := 0;
			else
				-- Holding two chips
				buffer_iq(pointer) <= chip_in;

				if pointer = 0 then
					pointer := pointer + 1;
					en_iq_out <= '0';
				elsif pointer = 1 then
					en_iq_out <= '1';
					pointer := 0;
				end if;
			end if;

		end if;
	end process;
	
	OUTPUT_SIGNALS: process(clk_1Mhz, en_iq_out, buffer_iq)
	begin
		if rising_edge(clk_1Mhz) then
			if reset = '1' then
				inphase <=  '0';
				quadrature <= '0';
			else
				-- Output signals for multiplication with sin,cos
				if en_iq_out = '1' then
				 	inphase <= buffer_iq(0);
				 	quadrature <= buffer_iq(1);
				end if;
			end if;
		end if;
	end process;
	
	--------------------------------------
	-- generation of a Tc delay
	--------------------------------------
	delay_buffer_chip(0) <= quadrature;

	gen_delay_en: for i in 1 to Delay generate
		delay_chip: process(clk_2Mhz)
			begin
				if rising_edge(clk_2Mhz) then
					delay_buffer_chip(i) <= delay_buffer_chip(i-1);
				end if;
			end process;
	end generate;

	quadrature_delayed <= delay_buffer_chip(Delay);

	--------------------------------------
	-- generation of sine&cos signals
	-- (not needed really - just for me)
	--------------------------------------
--	GEN_SINE: process(clk_sincos)
--		variable i : integer range 0 to 20 := 0;
--	begin
--		-- Each rise out a point of sine
--		if rising_edge(clk_sincos) then
--			if reset = '1' then
--				sine <= 0;
--				cos <= 0;
--				i := 0;
--			else
--				sine <= sine_values(i);
--				cos <= cos_values(i);
--				i := i + 1;
--				
--				if(i = 20) then
--					i := 0;
--				end if;
--			end if;
--		end if;
--	end process;

	--------------------------------------
	-- Multiplication of sine and chip
	-- Half-pulse shaping of chip data
	--------------------------------------
	MULT_CHIP_SIN: process(clk_sincos)
		variable j : integer range 0 to 20;
		variable w : integer range 0 to 20;
		variable h : integer range 0 to 20;
		variable y : integer range 0 to 20;
	begin
		-- Each rise, outputting a point of sine
		-- we output 20 values out of 21. 
		-- in sin it works due to the common point (0)
		-- but in cos we output 127, ..., 121. We are missing a value,
		-- we should output 127, ..., 127
		if rising_edge(clk_sincos) then
			if reset = '1' then
				modul_i <= 0;
				modul_q <= 0;
				j := 1;
				w := 10;
				h := 1;
				y := 10;
			else
				case inphase is
				   when '0' => 
					  -- ouputting 10 values.
					  -- 1-10 index
					  modul_i <= neg_sine_values(w);
					  if (w = 1) then
					      w := 10;
					  else
					      w := w - 1;
					  end if;

				   when others => 
					  -- ouputting 10 values.
					  -- 10-1 index
					  modul_i <= pos_sine_values(j);
					  if (j = 10) then
						  j := 1;
					  else
						  j := j + 1;
					  end if;
					  
			    end case;
	
				case quadrature_delayed is
				-- Look when signal changes state (1->0, 0->1)
				-- you have mistep, from 127 to -121 and from -127 to 121.
				-- because we dont have the commmon sample as in sin, the 0.
				   when '0' => 
					  -- Different LUT when signal is 0
					  modul_q <= neg_sine_values(y);
					  if (y = 1) then
					      y := 10;
					  else
					      y := y - 1;
					  end if;

				   when others => 
					  modul_q <= pos_sine_values(h);
					  if (h = 10) then
						  h := 1;
					  else
						  h := h + 1;
					  end if;
					  
			    end case;
				
		   end if;
				
		end if;
	end process;

	--------------------------------------
	-- Multiplication of sine and chip
	-- Half-pulse shaping of chip data
	--------------------------------------
	SUMMING_SIGNALS : process(clk_1Mhz)
	begin
		if rising_edge(clk_sincos) then
			if reset = '1' then
				sum <= 0;
			else
				sum <= modul_i + modul_q;
			end if;
		end if;
	end process;

end Behavioral;

